library verilog;
use verilog.vl_types.all;
entity memoria_vlg_check_tst is
    port(
        out0            : in     vl_logic;
        out1            : in     vl_logic;
        out2            : in     vl_logic;
        out3            : in     vl_logic;
        out4            : in     vl_logic;
        out5            : in     vl_logic;
        out6            : in     vl_logic;
        out7            : in     vl_logic;
        out8            : in     vl_logic;
        out9            : in     vl_logic;
        out10           : in     vl_logic;
        out11           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end memoria_vlg_check_tst;
