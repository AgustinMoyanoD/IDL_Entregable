library verilog;
use verilog.vl_types.all;
entity SumadorReCompleto123 is
    port(
        S_src0          : out    vl_logic;
        M0              : in     vl_logic;
        b0              : in     vl_logic;
        S_src1          : out    vl_logic;
        M1              : in     vl_logic;
        S_src2          : out    vl_logic;
        M2              : in     vl_logic;
        b2              : in     vl_logic;
        S_src3          : out    vl_logic;
        M3              : in     vl_logic;
        S_src4          : out    vl_logic;
        M4              : in     vl_logic;
        S_src5          : out    vl_logic;
        M5              : in     vl_logic;
        S_src6          : out    vl_logic;
        M6              : in     vl_logic;
        S_src7          : out    vl_logic;
        M7              : in     vl_logic;
        S_src8          : out    vl_logic;
        M8              : in     vl_logic;
        S_src10         : out    vl_logic;
        M10             : in     vl_logic;
        M9              : in     vl_logic;
        S_src9          : out    vl_logic;
        S_src11         : out    vl_logic;
        M11             : in     vl_logic;
        S_src12         : out    vl_logic;
        b1              : in     vl_logic
    );
end SumadorReCompleto123;
