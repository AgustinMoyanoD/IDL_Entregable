library verilog;
use verilog.vl_types.all;
entity SumadorReCompleto123_vlg_check_tst is
    port(
        S_src0          : in     vl_logic;
        S_src1          : in     vl_logic;
        S_src2          : in     vl_logic;
        S_src3          : in     vl_logic;
        S_src4          : in     vl_logic;
        S_src5          : in     vl_logic;
        S_src6          : in     vl_logic;
        S_src7          : in     vl_logic;
        S_src8          : in     vl_logic;
        S_src9          : in     vl_logic;
        S_src10         : in     vl_logic;
        S_src11         : in     vl_logic;
        S_src12         : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end SumadorReCompleto123_vlg_check_tst;
