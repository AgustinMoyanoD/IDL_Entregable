library verilog;
use verilog.vl_types.all;
entity Incrementador_vlg_vec_tst is
end Incrementador_vlg_vec_tst;
