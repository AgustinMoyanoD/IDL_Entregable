library verilog;
use verilog.vl_types.all;
entity MaquinaControlMultiplex_vlg_vec_tst is
end MaquinaControlMultiplex_vlg_vec_tst;
