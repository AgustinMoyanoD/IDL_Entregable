library verilog;
use verilog.vl_types.all;
entity compa2bits_vlg_vec_tst is
end compa2bits_vlg_vec_tst;
