library verilog;
use verilog.vl_types.all;
entity ffdConEnable_vlg_vec_tst is
end ffdConEnable_vlg_vec_tst;
