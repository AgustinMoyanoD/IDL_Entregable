library verilog;
use verilog.vl_types.all;
entity SemiSumador_vlg_check_tst is
    port(
        CryOut          : in     vl_logic;
        S               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end SemiSumador_vlg_check_tst;
