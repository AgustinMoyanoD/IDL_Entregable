library verilog;
use verilog.vl_types.all;
entity comparador12_vlg_vec_tst is
end comparador12_vlg_vec_tst;
