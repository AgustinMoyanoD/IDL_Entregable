library verilog;
use verilog.vl_types.all;
entity SemiSumador_vlg_vec_tst is
end SemiSumador_vlg_vec_tst;
