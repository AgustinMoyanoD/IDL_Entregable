library verilog;
use verilog.vl_types.all;
entity compa4bits_vlg_vec_tst is
end compa4bits_vlg_vec_tst;
