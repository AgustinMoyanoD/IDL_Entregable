library verilog;
use verilog.vl_types.all;
entity SumadorCompleto_vlg_check_tst is
    port(
        CryOut_sc       : in     vl_logic;
        S_sc            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end SumadorCompleto_vlg_check_tst;
