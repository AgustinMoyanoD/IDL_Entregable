library verilog;
use verilog.vl_types.all;
entity SumadorReCompleto123_vlg_vec_tst is
end SumadorReCompleto123_vlg_vec_tst;
