library verilog;
use verilog.vl_types.all;
entity SumadorReCompleto123_vlg_sample_tst is
    port(
        b0              : in     vl_logic;
        b1              : in     vl_logic;
        b2              : in     vl_logic;
        M0              : in     vl_logic;
        M1              : in     vl_logic;
        M2              : in     vl_logic;
        M3              : in     vl_logic;
        M4              : in     vl_logic;
        M5              : in     vl_logic;
        M6              : in     vl_logic;
        M7              : in     vl_logic;
        M8              : in     vl_logic;
        M9              : in     vl_logic;
        M10             : in     vl_logic;
        M11             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end SumadorReCompleto123_vlg_sample_tst;
