library verilog;
use verilog.vl_types.all;
entity memoria is
    port(
        out11           : out    vl_logic;
        CLK             : in     vl_logic;
        in11            : in     vl_logic;
        out10           : out    vl_logic;
        in10            : in     vl_logic;
        out9            : out    vl_logic;
        in9             : in     vl_logic;
        out8            : out    vl_logic;
        in8             : in     vl_logic;
        out7            : out    vl_logic;
        in7             : in     vl_logic;
        out6            : out    vl_logic;
        in6             : in     vl_logic;
        out5            : out    vl_logic;
        in5             : in     vl_logic;
        out4            : out    vl_logic;
        in4             : in     vl_logic;
        out3            : out    vl_logic;
        in3             : in     vl_logic;
        out2            : out    vl_logic;
        in2             : in     vl_logic;
        out1            : out    vl_logic;
        in1             : in     vl_logic;
        out0            : out    vl_logic;
        in0             : in     vl_logic
    );
end memoria;
