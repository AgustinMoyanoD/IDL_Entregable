library verilog;
use verilog.vl_types.all;
entity Cargador_vlg_check_tst is
    port(
        vf0             : in     vl_logic;
        vf1             : in     vl_logic;
        vf2             : in     vl_logic;
        vf3             : in     vl_logic;
        vf4             : in     vl_logic;
        vf5             : in     vl_logic;
        vf6             : in     vl_logic;
        vf7             : in     vl_logic;
        vf8             : in     vl_logic;
        vf9             : in     vl_logic;
        vf10            : in     vl_logic;
        vf11            : in     vl_logic;
        vi0             : in     vl_logic;
        vi1             : in     vl_logic;
        vi2             : in     vl_logic;
        vi3             : in     vl_logic;
        vi4             : in     vl_logic;
        vi5             : in     vl_logic;
        vi6             : in     vl_logic;
        vi7             : in     vl_logic;
        vi8             : in     vl_logic;
        vi9             : in     vl_logic;
        vi10            : in     vl_logic;
        vi11            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Cargador_vlg_check_tst;
