library verilog;
use verilog.vl_types.all;
entity compa8bits_vlg_vec_tst is
end compa8bits_vlg_vec_tst;
