library verilog;
use verilog.vl_types.all;
entity Cargador_vlg_vec_tst is
end Cargador_vlg_vec_tst;
